module main (CH, clock, reset, hsync, vsync, red, green, blue, sync, clk, blank);
	input [9:0] CH;
	input clock;
	input reset;
	output wire hsync;
	output wire vsync;
	output [7:0] red;
	output [7:0] green;
	output [7:0] blue;
	output sync;
	output clk;
	output blank;
	
	wire [7:0] color;
	assign color[0] = CH[0];
	assign color[1] = CH[1];
	assign color[2] = CH[2];
	assign color[3] = CH[3];
	assign color[4] = CH[4];
	assign color[5] = CH[5];
	assign color[6] = CH[6];
	assign color[7] = CH[7];
	
	clkdivider1 (clock, 0, clk25);
	
	ModuloVgaRoteiro (
		.clock(clock),
		.reset(!reset),
		.color_in(color),
		.next_x(),
		.next_y(),
		.hsync(hsync),
		.vsync(vsync),
		.red(red),
		.green(green),
		.blue(blue),
		.sync(sync),
		.clk(clk25),
		.blank(blank)
	);
endmodule